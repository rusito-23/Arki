module imem #(parameter N = 64)
				(input logic [5:0] addr, output logic [N-1:0] q);

endmodule
