
/**
* Execute Stage:
* Runs the given instruction (after being decoded).
*/

module execute(input logic ALUSrc,
					input logic [3:0] ALUControl,
					input logic [63:0] PC_E,
					input logic [63:0] signImm_E,
					input logic [63:0] readData1_E,
					input logic [63:0] readData2_E,
					output logic [63:0] PCBranch_E,
					output logic [63:0] aluResult_E,
					output logic [63:0] writeData_E,
					output logic zero_E)
					
	

endmodule
