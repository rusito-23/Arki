
module fetch(input logic PCSrc_F,
				 input logic clk,
				 input logic reset,
				 input logic [63:0] PCBranch_F,
				 output logic [63:0] imem_addr_F);
				 
	
				 
endmodule
